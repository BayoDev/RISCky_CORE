
module RV32_core(
    input clk
);

// wire we;
// reg [31:0] a,b;

// RAM ram_values(we,clk,a,b);

endmodule