

module top_bench
#(
    parameter XLEN = 32
)
(
	input                        in_clk,
    input                        rst,
	input                        uart_rx,
	output                       uart_tx,

    output leddington
);

reg [23:0] counter;

// Counter width calculation:
// 2^24 = 16,777,216 > 13,500,000
// So 24 bits is sufficient

always @(posedge in_clk or negedge rst) begin
    if (!rst) begin
        counter <= 24'd0;
        clk <= 1'b0;
    end
    else begin
        if (counter == 24'd13_499_999) begin
            counter <= 24'd0;
            clk <= ~clk;  // Toggle the output clock
        end
        else begin
            counter <= counter + 24'd1;
        end
    end
end

// reg clk,rst;
// always #5 clk = ~clk; 

// assign leddington = rst;
// assign leddington = tx_data[0];
assign leddington = clk;

integer i;

// COPIED DATA

parameter                        CLK_FRE  = 27;//Mhz
parameter                        UART_FRE = 115200;//Mhz
wire rx_data_ready = 1'b1;//always can receive data,
wire tx_data_ready;

// wire [7:0] rx_data;
// wire rx_data_valid;

// uart_rx#
// (
// 	.CLK_FRE(CLK_FRE),
// 	.BAUD_RATE(UART_FRE)
// ) uart_rx_inst
// (
// 	.clk                        (clk                      ),
// 	.rst_n                      (rst                      ),
// 	.rx_data                    (rx_data                  ),
// 	.rx_data_valid              (rx_data_valid            ),
// 	.rx_data_ready              (rx_data_ready            ),
// 	.rx_pin                     (uart_rx                  )
// );

wire tx_data_valid;
wire [7:0] tx_data;

uart_tx#
(
	.CLK_FRE(CLK_FRE),
	.BAUD_RATE(UART_FRE)
) uart_tx_inst
(
	.clk                        (clk                      ),
	.rst_n                      (rst                      ),
	.tx_data                    (tx_data                  ),
	.tx_data_valid              (tx_data_valid            ),
	.tx_data_ready              (tx_data_ready            ),
	.tx_pin                     (uart_tx                  )
);

// ==========================

//=======================
//      STAGE WIRES
//=======================

// IF

// input
wire [XLEN-1:0] if_branch_result_in;
wire if_was_branch_in;

// output
wire [31:0] if_instr_out;
wire [XLEN-1:0] if_pc_propagation_out;

// ID

// input
wire [31:0]     id_instr_in;
wire [4:0]      id_write_reg_dest_in;
wire            id_write_en_in;
wire [XLEN-1:0]     id_write_value_in;
wire [XLEN-1:0]     id_pc_propagation_in;

// output
wire [XLEN-1:0]     id_first_reg_out;
wire [XLEN-1:0]     id_second_reg_out;
wire [4:0]      id_write_reg_dest_out;
wire            id_write_en_out;
wire            id_reg_write_from_load;
wire [XLEN-1:0]     id_pc_propagation_out;
wire [2:0]      id_alu_op_base_out;
wire [6:0]      id_alu_op_ext_out;
wire            id_alu_src_out;
wire            id_is_branch_out;
wire            id_is_write_back;
wire            id_mem_write_out;
wire            id_mem_read_out;
wire [XLEN-1:0]     id_imm_value_out;
wire [2:0]   id_funct3_prop_out;
wire                id_is_link_and_jump_out;
wire                id_is_link_and_jump_reg_out;
wire                id_is_lui_out;
wire                id_is_auipc_out;

// EX

// input
wire [XLEN-1:0]     ex_op1_in;
wire [XLEN-1:0]     ex_op2_in;
wire [XLEN-1:0]     ex_sign_extended_in;
wire [2:0]      ex_alu_op_base_in;
wire [6:0]      ex_alu_op_ext_in;
wire            ex_alu_src_in;
wire [XLEN-1:0]     ex_pc_propagation_in;
wire            ex_is_branch_in;
wire [XLEN-1:0]     ex_imm_value_in;
wire [2:0]          ex_funct3_prop_in;
wire                ex_is_link_and_jump_in;
wire                ex_is_link_and_jump_reg_in;
wire                ex_is_lui_in;
wire                ex_is_auipc_in;

// output
wire [XLEN-1:0]     ex_result_out;
wire            ex_zero_out;
wire [XLEN-1:0]     ex_branch_result_out;
wire [XLEN-1:0]     ex_second_reg_propagation_out;
wire            ex_is_branch_out;
wire [2:0]      ex_funct3_prop_out;

// MEM

// input

wire [XLEN-1:0]     mem_ex_result_in;
wire            mem_ex_zero_in;
wire            mem_is_branch_op_in;
wire            mem_is_mem_write_in;
wire            mem_is_mem_read_in;
wire [XLEN-1:0]     mem_write_data_in;
wire            mem_dest_reg_prog_in;
wire [2:0]      mem_funct3_prop_in;

// output
wire            mem_is_valid_branch_out;
wire            mem_dest_reg_prog_out;
wire [XLEN-1:0]     mem_memory_res_out;
wire [XLEN-1:0]     mem_original_value_out;

// WB 

// input
wire            wb_mem_to_reg_in;
wire [XLEN-1:0]     wb_data_in;
wire [XLEN-1:0]     wb_orig_in;

// output
wire [XLEN-1:0]     wb_result_out;

instruction_fetch 
#(
    .XLEN(XLEN)
)
if_phase(
    .clk(clk),
    .rst(rst),

    .branch_result(if_branch_result_in),
    .was_branch(if_was_branch_in),

    .instr_out(if_instr_out),
    .pc_propagation(if_pc_propagation_out)
);

assign id_instr_in = if_instr_out;
assign id_pc_propagation_in = if_pc_propagation_out;

instruction_decoding 
#(
    .XLEN(XLEN)
)
id_phase(
    .clk(clk),
    .rst(rst),
    
    .instruction(id_instr_in),
    .reg_write_dest(id_write_reg_dest_in),
    .need_to_write(id_write_en_in),
    .reg_write_dest_value(id_write_value_in),

    .in_pc_value(id_pc_propagation_in),

    .first_reg(id_first_reg_out),
    .second_reg(id_second_reg_out),
    
    .reg_write_target(id_write_reg_dest_out),
    .reg_write(id_write_en_out),
    .reg_write_from_load(id_reg_write_from_load),

    .out_pc_value(id_pc_propagation_out),
    .ALU_op_base(id_alu_op_base_out),
    .ALU_op_ext(id_alu_op_ext_out),
    .ALU_src(id_alu_src_out),
    .imm_value(id_imm_value_out),

    .is_branch(id_is_branch_out),
    .mem_write(id_mem_write_out),
    .mem_read(id_mem_read_out),
    .is_write_back(id_is_write_back),

    .funct3_prop_out(id_funct3_prop_out),
    .is_link_and_jump(id_is_link_and_jump_out),
    .is_link_and_jump_reg(id_is_link_and_jump_reg_out),

    .is_lui(id_is_lui_out),
    .is_auipc(id_is_auipc_out)
);
// TODO: this is very messed up, this should be propagated through the ex phase
assign id_write_reg_dest_in = id_write_reg_dest_out;

assign ex_op1_in = id_first_reg_out;
assign ex_op2_in = id_second_reg_out;
assign ex_alu_src_in = id_alu_src_out;
assign ex_alu_op_base_in = id_alu_op_base_out;
assign ex_alu_op_ext_in = id_alu_op_ext_out;
assign ex_pc_propagation_in = id_pc_propagation_out;
assign ex_is_branch_in = id_is_branch_out;
assign ex_imm_value_in = id_imm_value_out;
assign ex_funct3_prop_in = id_funct3_prop_out;
assign ex_is_link_and_jump_in = id_is_link_and_jump_out;
assign ex_is_link_and_jump_reg_in = id_is_link_and_jump_reg_out;
assign ex_is_lui_in = id_is_lui_out;
assign ex_is_auipc_in = id_is_auipc_out;


execution 
#(
    .XLEN(XLEN)
)
ex_phase(
    .clk(clk),
    .rst(rst),

    .op1(ex_op1_in),
    .op2(ex_op2_in),

    .ALU_op(ex_alu_op_base_in),
    .ALU_op_ext(ex_alu_op_ext_in),
    .ALU_src(ex_alu_src_in),
    .imm_value(ex_imm_value_in),

    .funct3_prop_in(ex_funct3_prop_in),

    .is_link_and_jump(ex_is_link_and_jump_in),
    .is_link_and_jump_reg(ex_is_link_and_jump_reg_in),

    .is_lui(ex_is_lui_in),
    .is_auipc(ex_is_auipc_in),

    .res(ex_result_out),
    .zero(ex_zero_out),

    .in_pc_value(ex_pc_propagation_in),
    .is_branch_in(ex_is_branch_in),

    .branch_result(ex_branch_result_out),
    .second_reg_propagation(ex_second_reg_propagation_out),
    .is_branch_out(ex_is_branch_out),

    .funct3_prop_out(ex_funct3_prop_out)
);
// TODO: change this to go through mem for pipelining
assign if_branch_result_in = ex_branch_result_out;

assign mem_ex_result_in = ex_result_out;
assign mem_ex_zero_in = ex_zero_out;
assign mem_write_data_in = ex_second_reg_propagation_out;
assign if_was_branch_in = ex_is_branch_out;
assign mem_is_mem_write_in = id_mem_write_out;
assign mem_is_mem_read_in = id_mem_read_out;
assign mem_is_branch_op_in = id_is_branch_out;
assign mem_funct3_prop_in = ex_funct3_prop_out;

memory_access
#(
    .XLEN(XLEN)
)
mem_phase(
    .clk(clk),
    .rst(rst),

    .ex_result(mem_ex_result_in),
    .ex_zero(mem_ex_zero_in),
    .is_branch_op(mem_is_branch_op_in),
    .mem_write(mem_is_mem_write_in),
    .mem_read(mem_is_mem_read_in),
    .write_data(mem_write_data_in),
    .dest_reg_prog_in(mem_dest_reg_prog_in),

    .funct3_prop_in(mem_funct3_prop_in),

    .is_valid_branch(mem_is_valid_branch_out),
    .dest_reg_prog_out(mem_dest_reg_prog_out),
    .memory_res(mem_memory_res_out),
    .original_value(mem_original_value_out),

    .uart_tx_out(tx_data),
    .uart_tx_ready(tx_data_valid),

    .is_special(leddington2)
);
// TODO: change this to go through barrier with pipeline
// assign id_write_reg_dest_in = mem_dest_reg_prog_out;
assign id_write_en_in = id_write_en_out;

// assign wb_mem_to_reg_in 
assign wb_mem_to_reg_in = id_reg_write_from_load;
assign wb_data_in = mem_memory_res_out;
assign wb_orig_in = mem_original_value_out;
assign id_write_value_in = wb_result_out;

write_back
#(
    .XLEN(XLEN)
)
wb_phase(
    .mem_to_reg(wb_mem_to_reg_in),
    .data(wb_data_in),
    .orig(wb_orig_in),

    .result(wb_result_out)
);

// initial begin
//     $dumpfile("test.vcd");
//     $dumpvars(0,top_bench);

//     clk = 0;
//     rst=0;
//     #1 rst = 1;
//     #10 rst = 0;
//     #1000 $finish;
// end

endmodule