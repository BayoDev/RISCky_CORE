
module write_back(

    input mem_to_reg,

    
);



endmodule