
module memory_access(

    input clk,rst,

    input [31:0]    ex_result,
    input           ex_zero,
    input           mem_read,
    input           mem_write

    // output [31:0]   

);

// data_memory mem(

//     .clk(clk),
//     .rst(rst),

//     .address(),
//     .data_out()

// );



endmodule